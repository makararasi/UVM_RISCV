// TODO : add licence in all files

package test_pkg;
    import uvm_pkg::*;
    import seq_pkg::*;
    import riscv_mem_pkg::*;
    `include "uvm_macros.svh"

    `include "env.svh"
    `include "test_base.svh"

endpackage
