typedef uvm_sequencer #(riscv_seq_item) riscv_seqr;
