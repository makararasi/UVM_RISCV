// TODO : add licence in all files

package riscv_mem_pkg;
    import uvm_pkg::*;
    import seq_pkg::*;
    `include "uvm_macros.svh"
    `include "riscv_mem_driver.svh"
    `include "riscv_mem_monitor.svh"
    `include "riscv_mem_agent.svh"

endpackage

`include "riscv_mem_if.sv"
